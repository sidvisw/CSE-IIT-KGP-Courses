`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.11.2022 12:25:19
// Design Name: 
// Module Name: control_fsm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control_fsm(input clk, input rst, input indicator, input[31:0] x_comp, input[7:0] add_out, input cout, output reg[7:0] add_1, output reg[7:0] add_2, output reg cin,output reg en);

reg[11:0] pstate,nstate;

always@(posedge clk)
    begin
        if(rst)
            pstate<=6'd0;
        else
            pstate<=nstate;
    end

always@(*)
    begin
        case(pstate)
        12'd0:nstate<=12'd1;
        12'd1:nstate<=12'd2;
        12'd2:nstate<=12'd3;
        12'd3:nstate<=12'd4;
        12'd4:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd5;
                end
        12'd5:nstate<=12'd6;
        12'd6:nstate<=12'd7;
        12'd7:nstate<=12'd8;
        12'd8:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd9;
                end
        12'd9:nstate<=12'd10;
        12'd10:nstate<=12'd11;
        12'd11:nstate<=12'd12;
        12'd12:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd13;
                end
        12'd13:nstate<=12'd14;
        12'd14:nstate<=12'd15;
        12'd15:nstate<=12'd16;
        12'd16:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd17;
                end
        12'd17:nstate<=12'd18;
        12'd18:nstate<=12'd19;
        12'd19:nstate<=12'd20;
        12'd20:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd21;
                end
        12'd21:nstate<=12'd22;
        12'd22:nstate<=12'd23;
        12'd23:nstate<=12'd24;
        12'd24:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd25;
                end
        12'd25:nstate<=12'd26;
        12'd26:nstate<=12'd27;
        12'd27:nstate<=12'd28;
        12'd28:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd29;
                end
        12'd29:nstate<=12'd30;
        12'd30:nstate<=12'd31;
        12'd31:nstate<=12'd32;
        12'd32:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd33;
                end
        12'd33:nstate<=12'd34;
        12'd34:nstate<=12'd35;
        12'd35:nstate<=12'd36;
        12'd36:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd37;
                end
        12'd37:nstate<=12'd38;
        12'd38:nstate<=12'd39;
        12'd39:nstate<=12'd40;
        12'd40:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd41;
                end
        12'd41:nstate<=12'd42;
        12'd42:nstate<=12'd43;
        12'd43:nstate<=12'd44;
        12'd44:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd45;
                end
        12'd45:nstate<=12'd46;
        12'd46:nstate<=12'd47;
        12'd47:nstate<=12'd48;
        12'd48:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd49;
                end
        12'd49:nstate<=12'd50;
        12'd50:nstate<=12'd51;
        12'd51:nstate<=12'd52;
        12'd52:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd53;
                end
        12'd53:nstate<=12'd54;
        12'd54:nstate<=12'd55;
        12'd55:nstate<=12'd56;
        12'd56:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd57;
                end
        12'd57:nstate<=12'd58;
        12'd58:nstate<=12'd59;
        12'd59:nstate<=12'd60;
        12'd60:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd61;
                end
        12'd61:nstate<=12'd62;
        12'd62:nstate<=12'd63;
        12'd63:nstate<=12'd64;
        12'd64:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd65;
                end
        12'd65:nstate<=12'd66;
        12'd66:nstate<=12'd67;
        12'd67:nstate<=12'd68;
        12'd68:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd69;
                end
        12'd69:nstate<=12'd70;
        12'd70:nstate<=12'd71;
        12'd71:nstate<=12'd72;
        12'd72:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd73;
                end
        12'd73:nstate<=12'd74;
        12'd74:nstate<=12'd75;
        12'd75:nstate<=12'd76;
        12'd76:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd77;
                end
        12'd77:nstate<=12'd78;
        12'd78:nstate<=12'd79;
        12'd79:nstate<=12'd80;
        12'd80:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd81;
                end
        12'd81:nstate<=12'd82;
        12'd82:nstate<=12'd83;
        12'd83:nstate<=12'd84;
        12'd84:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd85;
                end
        12'd85:nstate<=12'd86;
        12'd86:nstate<=12'd87;
        12'd87:nstate<=12'd88;
        12'd88:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd89;
                end
        12'd89:nstate<=12'd90;
        12'd90:nstate<=12'd91;
        12'd91:nstate<=12'd92;
        12'd92:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd93;
                end
        12'd93:nstate<=12'd94;
        12'd94:nstate<=12'd95;
        12'd95:nstate<=12'd96;
        12'd96:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd97;
                end
        12'd97:nstate<=12'd98;
        12'd98:nstate<=12'd99;
        12'd99:nstate<=12'd100;
        12'd100:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd101;
                end
        12'd101:nstate<=12'd102;
        12'd102:nstate<=12'd103;
        12'd103:nstate<=12'd104;
        12'd104:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd105;
                end
        12'd105:nstate<=12'd106;
        12'd106:nstate<=12'd107;
        12'd107:nstate<=12'd108;
        12'd108:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd109;
                end
        12'd109:nstate<=12'd110;
        12'd110:nstate<=12'd111;
        12'd111:nstate<=12'd112;
        12'd112:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd113;
                end
        12'd113:nstate<=12'd114;
        12'd114:nstate<=12'd115;
        12'd115:nstate<=12'd116;
        12'd116:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd117;
                end
        12'd117:nstate<=12'd118;
        12'd118:nstate<=12'd119;
        12'd119:nstate<=12'd120;
        12'd120:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd121;
                end
        12'd121:nstate<=12'd122;
        12'd122:nstate<=12'd123;
        12'd123:nstate<=12'd124;
        12'd124:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd125;
                end
        12'd125:nstate<=12'd126;
        12'd126:nstate<=12'd127;
        12'd127:nstate<=12'd128;
        12'd128:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd129;
                end
        12'd129:nstate<=12'd130;
        12'd130:nstate<=12'd131;
        12'd131:nstate<=12'd132;
        12'd132:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd133;
                end
        12'd133:nstate<=12'd134;
        12'd134:nstate<=12'd135;
        12'd135:nstate<=12'd136;
        12'd136:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd137;
                end
        12'd137:nstate<=12'd138;
        12'd138:nstate<=12'd139;
        12'd139:nstate<=12'd140;
        12'd140:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd141;
                end
        12'd141:nstate<=12'd142;
        12'd142:nstate<=12'd143;
        12'd143:nstate<=12'd144;
        12'd144:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd145;
                end
        12'd145:nstate<=12'd146;
        12'd146:nstate<=12'd147;
        12'd147:nstate<=12'd148;
        12'd148:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd149;
                end
        12'd149:nstate<=12'd150;
        12'd150:nstate<=12'd151;
        12'd151:nstate<=12'd152;
        12'd152:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd153;
                end
        12'd153:nstate<=12'd154;
        12'd154:nstate<=12'd155;
        12'd155:nstate<=12'd156;
        12'd156:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd157;
                end
        12'd157:nstate<=12'd158;
        12'd158:nstate<=12'd159;
        12'd159:nstate<=12'd160;
        12'd160:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd161;
                end
        12'd161:nstate<=12'd162;
        12'd162:nstate<=12'd163;
        12'd163:nstate<=12'd164;
        12'd164:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd165;
                end
        12'd165:nstate<=12'd166;
        12'd166:nstate<=12'd167;
        12'd167:nstate<=12'd168;
        12'd168:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd169;
                end
        12'd169:nstate<=12'd170;
        12'd170:nstate<=12'd171;
        12'd171:nstate<=12'd172;
        12'd172:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd173;
                end
        12'd173:nstate<=12'd174;
        12'd174:nstate<=12'd175;
        12'd175:nstate<=12'd176;
        12'd176:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd177;
                end
        12'd177:nstate<=12'd178;
        12'd178:nstate<=12'd179;
        12'd179:nstate<=12'd180;
        12'd180:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd181;
                end
        12'd181:nstate<=12'd182;
        12'd182:nstate<=12'd183;
        12'd183:nstate<=12'd184;
        12'd184:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd185;
                end
        12'd185:nstate<=12'd186;
        12'd186:nstate<=12'd187;
        12'd187:nstate<=12'd188;
        12'd188:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd189;
                end
        12'd189:nstate<=12'd190;
        12'd190:nstate<=12'd191;
        12'd191:nstate<=12'd192;
        12'd192:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd193;
                end
        12'd193:nstate<=12'd194;
        12'd194:nstate<=12'd195;
        12'd195:nstate<=12'd196;
        12'd196:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd197;
                end
        12'd197:nstate<=12'd198;
        12'd198:nstate<=12'd199;
        12'd199:nstate<=12'd200;
        12'd200:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd201;
                end
        12'd201:nstate<=12'd202;
        12'd202:nstate<=12'd203;
        12'd203:nstate<=12'd204;
        12'd204:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd205;
                end
        12'd205:nstate<=12'd206;
        12'd206:nstate<=12'd207;
        12'd207:nstate<=12'd208;
        12'd208:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd209;
                end
        12'd209:nstate<=12'd210;
        12'd210:nstate<=12'd211;
        12'd211:nstate<=12'd212;
        12'd212:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd213;
                end
        12'd213:nstate<=12'd214;
        12'd214:nstate<=12'd215;
        12'd215:nstate<=12'd216;
        12'd216:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd217;
                end
        12'd217:nstate<=12'd218;
        12'd218:nstate<=12'd219;
        12'd219:nstate<=12'd220;
        12'd220:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd221;
                end
        12'd221:nstate<=12'd222;
        12'd222:nstate<=12'd223;
        12'd223:nstate<=12'd224;
        12'd224:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd225;
                end
        12'd225:nstate<=12'd226;
        12'd226:nstate<=12'd227;
        12'd227:nstate<=12'd228;
        12'd228:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd229;
                end
        12'd229:nstate<=12'd230;
        12'd230:nstate<=12'd231;
        12'd231:nstate<=12'd232;
        12'd232:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd233;
                end
        12'd233:nstate<=12'd234;
        12'd234:nstate<=12'd235;
        12'd235:nstate<=12'd236;
        12'd236:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd237;
                end
        12'd237:nstate<=12'd238;
        12'd238:nstate<=12'd239;
        12'd239:nstate<=12'd240;
        12'd240:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd241;
                end
        12'd241:nstate<=12'd242;
        12'd242:nstate<=12'd243;
        12'd243:nstate<=12'd244;
        12'd244:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd245;
                end
        12'd245:nstate<=12'd246;
        12'd246:nstate<=12'd247;
        12'd247:nstate<=12'd248;
        12'd248:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd249;
                end
        12'd249:nstate<=12'd250;
        12'd250:nstate<=12'd251;
        12'd251:nstate<=12'd252;
        12'd252:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd253;
                end
        12'd253:nstate<=12'd254;
        12'd254:nstate<=12'd255;
        12'd255:nstate<=12'd256;
        12'd256:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd257;
                end
        12'd257:nstate<=12'd258;
        12'd258:nstate<=12'd259;
        12'd259:nstate<=12'd260;
        12'd260:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd261;
                end
        12'd261:nstate<=12'd262;
        12'd262:nstate<=12'd263;
        12'd263:nstate<=12'd264;
        12'd264:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd265;
                end
        12'd265:nstate<=12'd266;
        12'd266:nstate<=12'd267;
        12'd267:nstate<=12'd268;
        12'd268:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd269;
                end
        12'd269:nstate<=12'd270;
        12'd270:nstate<=12'd271;
        12'd271:nstate<=12'd272;
        12'd272:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd273;
                end
        12'd273:nstate<=12'd274;
        12'd274:nstate<=12'd275;
        12'd275:nstate<=12'd276;
        12'd276:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd277;
                end
        12'd277:nstate<=12'd278;
        12'd278:nstate<=12'd279;
        12'd279:nstate<=12'd280;
        12'd280:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd281;
                end
        12'd281:nstate<=12'd282;
        12'd282:nstate<=12'd283;
        12'd283:nstate<=12'd284;
        12'd284:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd285;
                end
        12'd285:nstate<=12'd286;
        12'd286:nstate<=12'd287;
        12'd287:nstate<=12'd288;
        12'd288:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd289;
                end
        12'd289:nstate<=12'd290;
        12'd290:nstate<=12'd291;
        12'd291:nstate<=12'd292;
        12'd292:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd293;
                end
        12'd293:nstate<=12'd294;
        12'd294:nstate<=12'd295;
        12'd295:nstate<=12'd296;
        12'd296:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd297;
                end
        12'd297:nstate<=12'd298;
        12'd298:nstate<=12'd299;
        12'd299:nstate<=12'd300;
        12'd300:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd301;
                end
        12'd301:nstate<=12'd302;
        12'd302:nstate<=12'd303;
        12'd303:nstate<=12'd304;
        12'd304:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd305;
                end
        12'd305:nstate<=12'd306;
        12'd306:nstate<=12'd307;
        12'd307:nstate<=12'd308;
        12'd308:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd309;
                end
        12'd309:nstate<=12'd310;
        12'd310:nstate<=12'd311;
        12'd311:nstate<=12'd312;
        12'd312:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd313;
                end
        12'd313:nstate<=12'd314;
        12'd314:nstate<=12'd315;
        12'd315:nstate<=12'd316;
        12'd316:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd317;
                end
        12'd317:nstate<=12'd318;
        12'd318:nstate<=12'd319;
        12'd319:nstate<=12'd320;
        12'd320:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd321;
                end
        12'd321:nstate<=12'd322;
        12'd322:nstate<=12'd323;
        12'd323:nstate<=12'd324;
        12'd324:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd325;
                end
        12'd325:nstate<=12'd326;
        12'd326:nstate<=12'd327;
        12'd327:nstate<=12'd328;
        12'd328:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd329;
                end
        12'd329:nstate<=12'd330;
        12'd330:nstate<=12'd331;
        12'd331:nstate<=12'd332;
        12'd332:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd333;
                end
        12'd333:nstate<=12'd334;
        12'd334:nstate<=12'd335;
        12'd335:nstate<=12'd336;
        12'd336:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd337;
                end
        12'd337:nstate<=12'd338;
        12'd338:nstate<=12'd339;
        12'd339:nstate<=12'd340;
        12'd340:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd341;
                end
        12'd341:nstate<=12'd342;
        12'd342:nstate<=12'd343;
        12'd343:nstate<=12'd344;
        12'd344:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd345;
                end
        12'd345:nstate<=12'd346;
        12'd346:nstate<=12'd347;
        12'd347:nstate<=12'd348;
        12'd348:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd349;
                end
        12'd349:nstate<=12'd350;
        12'd350:nstate<=12'd351;
        12'd351:nstate<=12'd352;
        12'd352:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd353;
                end
        12'd353:nstate<=12'd354;
        12'd354:nstate<=12'd355;
        12'd355:nstate<=12'd356;
        12'd356:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd357;
                end
        12'd357:nstate<=12'd358;
        12'd358:nstate<=12'd359;
        12'd359:nstate<=12'd360;
        12'd360:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd361;
                end
        12'd361:nstate<=12'd362;
        12'd362:nstate<=12'd363;
        12'd363:nstate<=12'd364;
        12'd364:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd365;
                end
        12'd365:nstate<=12'd366;
        12'd366:nstate<=12'd367;
        12'd367:nstate<=12'd368;
        12'd368:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd369;
                end
        12'd369:nstate<=12'd370;
        12'd370:nstate<=12'd371;
        12'd371:nstate<=12'd372;
        12'd372:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd373;
                end
        12'd373:nstate<=12'd374;
        12'd374:nstate<=12'd375;
        12'd375:nstate<=12'd376;
        12'd376:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd377;
                end
        12'd377:nstate<=12'd378;
        12'd378:nstate<=12'd379;
        12'd379:nstate<=12'd380;
        12'd380:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd381;
                end
        12'd381:nstate<=12'd382;
        12'd382:nstate<=12'd383;
        12'd383:nstate<=12'd384;
        12'd384:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd385;
                end
        12'd385:nstate<=12'd386;
        12'd386:nstate<=12'd387;
        12'd387:nstate<=12'd388;
        12'd388:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd389;
                end
        12'd389:nstate<=12'd390;
        12'd390:nstate<=12'd391;
        12'd391:nstate<=12'd392;
        12'd392:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd393;
                end
        12'd393:nstate<=12'd394;
        12'd394:nstate<=12'd395;
        12'd395:nstate<=12'd396;
        12'd396:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd397;
                end
        12'd397:nstate<=12'd398;
        12'd398:nstate<=12'd399;
        12'd399:nstate<=12'd400;
        12'd400:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd401;
                end
        12'd401:nstate<=12'd402;
        12'd402:nstate<=12'd403;
        12'd403:nstate<=12'd404;
        12'd404:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd405;
                end
        12'd405:nstate<=12'd406;
        12'd406:nstate<=12'd407;
        12'd407:nstate<=12'd408;
        12'd408:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd409;
                end
        12'd409:nstate<=12'd410;
        12'd410:nstate<=12'd411;
        12'd411:nstate<=12'd412;
        12'd412:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd413;
                end
        12'd413:nstate<=12'd414;
        12'd414:nstate<=12'd415;
        12'd415:nstate<=12'd416;
        12'd416:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd417;
                end
        12'd417:nstate<=12'd418;
        12'd418:nstate<=12'd419;
        12'd419:nstate<=12'd420;
        12'd420:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd421;
                end
        12'd421:nstate<=12'd422;
        12'd422:nstate<=12'd423;
        12'd423:nstate<=12'd424;
        12'd424:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd425;
                end
        12'd425:nstate<=12'd426;
        12'd426:nstate<=12'd427;
        12'd427:nstate<=12'd428;
        12'd428:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd429;
                end
        12'd429:nstate<=12'd430;
        12'd430:nstate<=12'd431;
        12'd431:nstate<=12'd432;
        12'd432:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd433;
                end
        12'd433:nstate<=12'd434;
        12'd434:nstate<=12'd435;
        12'd435:nstate<=12'd436;
        12'd436:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd437;
                end
        12'd437:nstate<=12'd438;
        12'd438:nstate<=12'd439;
        12'd439:nstate<=12'd440;
        12'd440:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd441;
                end
        12'd441:nstate<=12'd442;
        12'd442:nstate<=12'd443;
        12'd443:nstate<=12'd444;
        12'd444:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd445;
                end
        12'd445:nstate<=12'd446;
        12'd446:nstate<=12'd447;
        12'd447:nstate<=12'd448;
        12'd448:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd449;
                end
        12'd449:nstate<=12'd450;
        12'd450:nstate<=12'd451;
        12'd451:nstate<=12'd452;
        12'd452:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd453;
                end
        12'd453:nstate<=12'd454;
        12'd454:nstate<=12'd455;
        12'd455:nstate<=12'd456;
        12'd456:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd457;
                end
        12'd457:nstate<=12'd458;
        12'd458:nstate<=12'd459;
        12'd459:nstate<=12'd460;
        12'd460:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd461;
                end
        12'd461:nstate<=12'd462;
        12'd462:nstate<=12'd463;
        12'd463:nstate<=12'd464;
        12'd464:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd465;
                end
        12'd465:nstate<=12'd466;
        12'd466:nstate<=12'd467;
        12'd467:nstate<=12'd468;
        12'd468:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd469;
                end
        12'd469:nstate<=12'd470;
        12'd470:nstate<=12'd471;
        12'd471:nstate<=12'd472;
        12'd472:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd473;
                end
        12'd473:nstate<=12'd474;
        12'd474:nstate<=12'd475;
        12'd475:nstate<=12'd476;
        12'd476:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd477;
                end
        12'd477:nstate<=12'd478;
        12'd478:nstate<=12'd479;
        12'd479:nstate<=12'd480;
        12'd480:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd481;
                end
        12'd481:nstate<=12'd482;
        12'd482:nstate<=12'd483;
        12'd483:nstate<=12'd484;
        12'd484:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd485;
                end
        12'd485:nstate<=12'd486;
        12'd486:nstate<=12'd487;
        12'd487:nstate<=12'd488;
        12'd488:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd489;
                end
        12'd489:nstate<=12'd490;
        12'd490:nstate<=12'd491;
        12'd491:nstate<=12'd492;
        12'd492:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd493;
                end
        12'd493:nstate<=12'd494;
        12'd494:nstate<=12'd495;
        12'd495:nstate<=12'd496;
        12'd496:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd497;
                end
        12'd497:nstate<=12'd498;
        12'd498:nstate<=12'd499;
        12'd499:nstate<=12'd500;
        12'd500:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd501;
                end
        12'd501:nstate<=12'd502;
        12'd502:nstate<=12'd503;
        12'd503:nstate<=12'd504;
        12'd504:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd505;
                end
        12'd505:nstate<=12'd506;
        12'd506:nstate<=12'd507;
        12'd507:nstate<=12'd508;
        12'd508:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd509;
                end
        12'd509:nstate<=12'd510;
        12'd510:nstate<=12'd511;
        12'd511:nstate<=12'd512;
        12'd512:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd513;
                end
        12'd513:nstate<=12'd514;
        12'd514:nstate<=12'd515;
        12'd515:nstate<=12'd516;
        12'd516:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd517;
                end
        12'd517:nstate<=12'd518;
        12'd518:nstate<=12'd519;
        12'd519:nstate<=12'd520;
        12'd520:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd521;
                end
        12'd521:nstate<=12'd522;
        12'd522:nstate<=12'd523;
        12'd523:nstate<=12'd524;
        12'd524:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd525;
                end
        12'd525:nstate<=12'd526;
        12'd526:nstate<=12'd527;
        12'd527:nstate<=12'd528;
        12'd528:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd529;
                end
        12'd529:nstate<=12'd530;
        12'd530:nstate<=12'd531;
        12'd531:nstate<=12'd532;
        12'd532:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd533;
                end
        12'd533:nstate<=12'd534;
        12'd534:nstate<=12'd535;
        12'd535:nstate<=12'd536;
        12'd536:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd537;
                end
        12'd537:nstate<=12'd538;
        12'd538:nstate<=12'd539;
        12'd539:nstate<=12'd540;
        12'd540:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd541;
                end
        12'd541:nstate<=12'd542;
        12'd542:nstate<=12'd543;
        12'd543:nstate<=12'd544;
        12'd544:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd545;
                end
        12'd545:nstate<=12'd546;
        12'd546:nstate<=12'd547;
        12'd547:nstate<=12'd548;
        12'd548:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd549;
                end
        12'd549:nstate<=12'd550;
        12'd550:nstate<=12'd551;
        12'd551:nstate<=12'd552;
        12'd552:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd553;
                end
        12'd553:nstate<=12'd554;
        12'd554:nstate<=12'd555;
        12'd555:nstate<=12'd556;
        12'd556:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd557;
                end
        12'd557:nstate<=12'd558;
        12'd558:nstate<=12'd559;
        12'd559:nstate<=12'd560;
        12'd560:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd561;
                end
        12'd561:nstate<=12'd562;
        12'd562:nstate<=12'd563;
        12'd563:nstate<=12'd564;
        12'd564:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd565;
                end
        12'd565:nstate<=12'd566;
        12'd566:nstate<=12'd567;
        12'd567:nstate<=12'd568;
        12'd568:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd569;
                end
        12'd569:nstate<=12'd570;
        12'd570:nstate<=12'd571;
        12'd571:nstate<=12'd572;
        12'd572:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd573;
                end
        12'd573:nstate<=12'd574;
        12'd574:nstate<=12'd575;
        12'd575:nstate<=12'd576;
        12'd576:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd577;
                end
        12'd577:nstate<=12'd578;
        12'd578:nstate<=12'd579;
        12'd579:nstate<=12'd580;
        12'd580:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd581;
                end
        12'd581:nstate<=12'd582;
        12'd582:nstate<=12'd583;
        12'd583:nstate<=12'd584;
        12'd584:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd585;
                end
        12'd585:nstate<=12'd586;
        12'd586:nstate<=12'd587;
        12'd587:nstate<=12'd588;
        12'd588:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd589;
                end
        12'd589:nstate<=12'd590;
        12'd590:nstate<=12'd591;
        12'd591:nstate<=12'd592;
        12'd592:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd593;
                end
        12'd593:nstate<=12'd594;
        12'd594:nstate<=12'd595;
        12'd595:nstate<=12'd596;
        12'd596:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd597;
                end
        12'd597:nstate<=12'd598;
        12'd598:nstate<=12'd599;
        12'd599:nstate<=12'd600;
        12'd600:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd601;
                end
        12'd601:nstate<=12'd602;
        12'd602:nstate<=12'd603;
        12'd603:nstate<=12'd604;
        12'd604:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd605;
                end
        12'd605:nstate<=12'd606;
        12'd606:nstate<=12'd607;
        12'd607:nstate<=12'd608;
        12'd608:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd609;
                end
        12'd609:nstate<=12'd610;
        12'd610:nstate<=12'd611;
        12'd611:nstate<=12'd612;
        12'd612:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd613;
                end
        12'd613:nstate<=12'd614;
        12'd614:nstate<=12'd615;
        12'd615:nstate<=12'd616;
        12'd616:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd617;
                end
        12'd617:nstate<=12'd618;
        12'd618:nstate<=12'd619;
        12'd619:nstate<=12'd620;
        12'd620:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd621;
                end
        12'd621:nstate<=12'd622;
        12'd622:nstate<=12'd623;
        12'd623:nstate<=12'd624;
        12'd624:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd625;
                end
        12'd625:nstate<=12'd626;
        12'd626:nstate<=12'd627;
        12'd627:nstate<=12'd628;
        12'd628:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd629;
                end
        12'd629:nstate<=12'd630;
        12'd630:nstate<=12'd631;
        12'd631:nstate<=12'd632;
        12'd632:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd633;
                end
        12'd633:nstate<=12'd634;
        12'd634:nstate<=12'd635;
        12'd635:nstate<=12'd636;
        12'd636:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd637;
                end
        12'd637:nstate<=12'd638;
        12'd638:nstate<=12'd639;
        12'd639:nstate<=12'd640;
        12'd640:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd641;
                end
        12'd641:nstate<=12'd642;
        12'd642:nstate<=12'd643;
        12'd643:nstate<=12'd644;
        12'd644:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd645;
                end
        12'd645:nstate<=12'd646;
        12'd646:nstate<=12'd647;
        12'd647:nstate<=12'd648;
        12'd648:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd649;
                end
        12'd649:nstate<=12'd650;
        12'd650:nstate<=12'd651;
        12'd651:nstate<=12'd652;
        12'd652:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd653;
                end
        12'd653:nstate<=12'd654;
        12'd654:nstate<=12'd655;
        12'd655:nstate<=12'd656;
        12'd656:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd657;
                end
        12'd657:nstate<=12'd658;
        12'd658:nstate<=12'd659;
        12'd659:nstate<=12'd660;
        12'd660:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd661;
                end
        12'd661:nstate<=12'd662;
        12'd662:nstate<=12'd663;
        12'd663:nstate<=12'd664;
        12'd664:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd665;
                end
        12'd665:nstate<=12'd666;
        12'd666:nstate<=12'd667;
        12'd667:nstate<=12'd668;
        12'd668:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd669;
                end
        12'd669:nstate<=12'd670;
        12'd670:nstate<=12'd671;
        12'd671:nstate<=12'd672;
        12'd672:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd673;
                end
        12'd673:nstate<=12'd674;
        12'd674:nstate<=12'd675;
        12'd675:nstate<=12'd676;
        12'd676:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd677;
                end
        12'd677:nstate<=12'd678;
        12'd678:nstate<=12'd679;
        12'd679:nstate<=12'd680;
        12'd680:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd681;
                end
        12'd681:nstate<=12'd682;
        12'd682:nstate<=12'd683;
        12'd683:nstate<=12'd684;
        12'd684:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd685;
                end
        12'd685:nstate<=12'd686;
        12'd686:nstate<=12'd687;
        12'd687:nstate<=12'd688;
        12'd688:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd689;
                end
        12'd689:nstate<=12'd690;
        12'd690:nstate<=12'd691;
        12'd691:nstate<=12'd692;
        12'd692:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd693;
                end
        12'd693:nstate<=12'd694;
        12'd694:nstate<=12'd695;
        12'd695:nstate<=12'd696;
        12'd696:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd697;
                end
        12'd697:nstate<=12'd698;
        12'd698:nstate<=12'd699;
        12'd699:nstate<=12'd700;
        12'd700:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd701;
                end
        12'd701:nstate<=12'd702;
        12'd702:nstate<=12'd703;
        12'd703:nstate<=12'd704;
        12'd704:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd705;
                end
        12'd705:nstate<=12'd706;
        12'd706:nstate<=12'd707;
        12'd707:nstate<=12'd708;
        12'd708:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd709;
                end
        12'd709:nstate<=12'd710;
        12'd710:nstate<=12'd711;
        12'd711:nstate<=12'd712;
        12'd712:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd713;
                end
        12'd713:nstate<=12'd714;
        12'd714:nstate<=12'd715;
        12'd715:nstate<=12'd716;
        12'd716:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd717;
                end
        12'd717:nstate<=12'd718;
        12'd718:nstate<=12'd719;
        12'd719:nstate<=12'd720;
        12'd720:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd721;
                end
        12'd721:nstate<=12'd722;
        12'd722:nstate<=12'd723;
        12'd723:nstate<=12'd724;
        12'd724:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd725;
                end
        12'd725:nstate<=12'd726;
        12'd726:nstate<=12'd727;
        12'd727:nstate<=12'd728;
        12'd728:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd729;
                end
        12'd729:nstate<=12'd730;
        12'd730:nstate<=12'd731;
        12'd731:nstate<=12'd732;
        12'd732:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd733;
                end
        12'd733:nstate<=12'd734;
        12'd734:nstate<=12'd735;
        12'd735:nstate<=12'd736;
        12'd736:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd737;
                end
        12'd737:nstate<=12'd738;
        12'd738:nstate<=12'd739;
        12'd739:nstate<=12'd740;
        12'd740:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd741;
                end
        12'd741:nstate<=12'd742;
        12'd742:nstate<=12'd743;
        12'd743:nstate<=12'd744;
        12'd744:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd745;
                end
        12'd745:nstate<=12'd746;
        12'd746:nstate<=12'd747;
        12'd747:nstate<=12'd748;
        12'd748:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd749;
                end
        12'd749:nstate<=12'd750;
        12'd750:nstate<=12'd751;
        12'd751:nstate<=12'd752;
        12'd752:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd753;
                end
        12'd753:nstate<=12'd754;
        12'd754:nstate<=12'd755;
        12'd755:nstate<=12'd756;
        12'd756:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd757;
                end
        12'd757:nstate<=12'd758;
        12'd758:nstate<=12'd759;
        12'd759:nstate<=12'd760;
        12'd760:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd761;
                end
        12'd761:nstate<=12'd762;
        12'd762:nstate<=12'd763;
        12'd763:nstate<=12'd764;
        12'd764:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd765;
                end
        12'd765:nstate<=12'd766;
        12'd766:nstate<=12'd767;
        12'd767:nstate<=12'd768;
        12'd768:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd769;
                end
        12'd769:nstate<=12'd770;
        12'd770:nstate<=12'd771;
        12'd771:nstate<=12'd772;
        12'd772:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd773;
                end
        12'd773:nstate<=12'd774;
        12'd774:nstate<=12'd775;
        12'd775:nstate<=12'd776;
        12'd776:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd777;
                end
        12'd777:nstate<=12'd778;
        12'd778:nstate<=12'd779;
        12'd779:nstate<=12'd780;
        12'd780:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd781;
                end
        12'd781:nstate<=12'd782;
        12'd782:nstate<=12'd783;
        12'd783:nstate<=12'd784;
        12'd784:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd785;
                end
        12'd785:nstate<=12'd786;
        12'd786:nstate<=12'd787;
        12'd787:nstate<=12'd788;
        12'd788:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd789;
                end
        12'd789:nstate<=12'd790;
        12'd790:nstate<=12'd791;
        12'd791:nstate<=12'd792;
        12'd792:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd793;
                end
        12'd793:nstate<=12'd794;
        12'd794:nstate<=12'd795;
        12'd795:nstate<=12'd796;
        12'd796:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd797;
                end
        12'd797:nstate<=12'd798;
        12'd798:nstate<=12'd799;
        12'd799:nstate<=12'd800;
        12'd800:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd801;
                end
        12'd801:nstate<=12'd802;
        12'd802:nstate<=12'd803;
        12'd803:nstate<=12'd804;
        12'd804:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd805;
                end
        12'd805:nstate<=12'd806;
        12'd806:nstate<=12'd807;
        12'd807:nstate<=12'd808;
        12'd808:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd809;
                end
        12'd809:nstate<=12'd810;
        12'd810:nstate<=12'd811;
        12'd811:nstate<=12'd812;
        12'd812:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd813;
                end
        12'd813:nstate<=12'd814;
        12'd814:nstate<=12'd815;
        12'd815:nstate<=12'd816;
        12'd816:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd817;
                end
        12'd817:nstate<=12'd818;
        12'd818:nstate<=12'd819;
        12'd819:nstate<=12'd820;
        12'd820:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd821;
                end
        12'd821:nstate<=12'd822;
        12'd822:nstate<=12'd823;
        12'd823:nstate<=12'd824;
        12'd824:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd825;
                end
        12'd825:nstate<=12'd826;
        12'd826:nstate<=12'd827;
        12'd827:nstate<=12'd828;
        12'd828:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd829;
                end
        12'd829:nstate<=12'd830;
        12'd830:nstate<=12'd831;
        12'd831:nstate<=12'd832;
        12'd832:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd833;
                end
        12'd833:nstate<=12'd834;
        12'd834:nstate<=12'd835;
        12'd835:nstate<=12'd836;
        12'd836:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd837;
                end
        12'd837:nstate<=12'd838;
        12'd838:nstate<=12'd839;
        12'd839:nstate<=12'd840;
        12'd840:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd841;
                end
        12'd841:nstate<=12'd842;
        12'd842:nstate<=12'd843;
        12'd843:nstate<=12'd844;
        12'd844:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd845;
                end
        12'd845:nstate<=12'd846;
        12'd846:nstate<=12'd847;
        12'd847:nstate<=12'd848;
        12'd848:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd849;
                end
        12'd849:nstate<=12'd850;
        12'd850:nstate<=12'd851;
        12'd851:nstate<=12'd852;
        12'd852:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd853;
                end
        12'd853:nstate<=12'd854;
        12'd854:nstate<=12'd855;
        12'd855:nstate<=12'd856;
        12'd856:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd857;
                end
        12'd857:nstate<=12'd858;
        12'd858:nstate<=12'd859;
        12'd859:nstate<=12'd860;
        12'd860:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd861;
                end
        12'd861:nstate<=12'd862;
        12'd862:nstate<=12'd863;
        12'd863:nstate<=12'd864;
        12'd864:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd865;
                end
        12'd865:nstate<=12'd866;
        12'd866:nstate<=12'd867;
        12'd867:nstate<=12'd868;
        12'd868:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd869;
                end
        12'd869:nstate<=12'd870;
        12'd870:nstate<=12'd871;
        12'd871:nstate<=12'd872;
        12'd872:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd873;
                end
        12'd873:nstate<=12'd874;
        12'd874:nstate<=12'd875;
        12'd875:nstate<=12'd876;
        12'd876:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd877;
                end
        12'd877:nstate<=12'd878;
        12'd878:nstate<=12'd879;
        12'd879:nstate<=12'd880;
        12'd880:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd881;
                end
        12'd881:nstate<=12'd882;
        12'd882:nstate<=12'd883;
        12'd883:nstate<=12'd884;
        12'd884:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd885;
                end
        12'd885:nstate<=12'd886;
        12'd886:nstate<=12'd887;
        12'd887:nstate<=12'd888;
        12'd888:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd889;
                end
        12'd889:nstate<=12'd890;
        12'd890:nstate<=12'd891;
        12'd891:nstate<=12'd892;
        12'd892:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd893;
                end
        12'd893:nstate<=12'd894;
        12'd894:nstate<=12'd895;
        12'd895:nstate<=12'd896;
        12'd896:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd897;
                end
        12'd897:nstate<=12'd898;
        12'd898:nstate<=12'd899;
        12'd899:nstate<=12'd900;
        12'd900:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd901;
                end
        12'd901:nstate<=12'd902;
        12'd902:nstate<=12'd903;
        12'd903:nstate<=12'd904;
        12'd904:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd905;
                end
        12'd905:nstate<=12'd906;
        12'd906:nstate<=12'd907;
        12'd907:nstate<=12'd908;
        12'd908:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd909;
                end
        12'd909:nstate<=12'd910;
        12'd910:nstate<=12'd911;
        12'd911:nstate<=12'd912;
        12'd912:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd913;
                end
        12'd913:nstate<=12'd914;
        12'd914:nstate<=12'd915;
        12'd915:nstate<=12'd916;
        12'd916:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd917;
                end
        12'd917:nstate<=12'd918;
        12'd918:nstate<=12'd919;
        12'd919:nstate<=12'd920;
        12'd920:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd921;
                end
        12'd921:nstate<=12'd922;
        12'd922:nstate<=12'd923;
        12'd923:nstate<=12'd924;
        12'd924:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd925;
                end
        12'd925:nstate<=12'd926;
        12'd926:nstate<=12'd927;
        12'd927:nstate<=12'd928;
        12'd928:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd929;
                end
        12'd929:nstate<=12'd930;
        12'd930:nstate<=12'd931;
        12'd931:nstate<=12'd932;
        12'd932:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd933;
                end
        12'd933:nstate<=12'd934;
        12'd934:nstate<=12'd935;
        12'd935:nstate<=12'd936;
        12'd936:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd937;
                end
        12'd937:nstate<=12'd938;
        12'd938:nstate<=12'd939;
        12'd939:nstate<=12'd940;
        12'd940:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd941;
                end
        12'd941:nstate<=12'd942;
        12'd942:nstate<=12'd943;
        12'd943:nstate<=12'd944;
        12'd944:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd945;
                end
        12'd945:nstate<=12'd946;
        12'd946:nstate<=12'd947;
        12'd947:nstate<=12'd948;
        12'd948:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd949;
                end
        12'd949:nstate<=12'd950;
        12'd950:nstate<=12'd951;
        12'd951:nstate<=12'd952;
        12'd952:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd953;
                end
        12'd953:nstate<=12'd954;
        12'd954:nstate<=12'd955;
        12'd955:nstate<=12'd956;
        12'd956:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd957;
                end
        12'd957:nstate<=12'd958;
        12'd958:nstate<=12'd959;
        12'd959:nstate<=12'd960;
        12'd960:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd961;
                end
        12'd961:nstate<=12'd962;
        12'd962:nstate<=12'd963;
        12'd963:nstate<=12'd964;
        12'd964:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd965;
                end
        12'd965:nstate<=12'd966;
        12'd966:nstate<=12'd967;
        12'd967:nstate<=12'd968;
        12'd968:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd969;
                end
        12'd969:nstate<=12'd970;
        12'd970:nstate<=12'd971;
        12'd971:nstate<=12'd972;
        12'd972:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd973;
                end
        12'd973:nstate<=12'd974;
        12'd974:nstate<=12'd975;
        12'd975:nstate<=12'd976;
        12'd976:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd977;
                end
        12'd977:nstate<=12'd978;
        12'd978:nstate<=12'd979;
        12'd979:nstate<=12'd980;
        12'd980:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd981;
                end
        12'd981:nstate<=12'd982;
        12'd982:nstate<=12'd983;
        12'd983:nstate<=12'd984;
        12'd984:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd985;
                end
        12'd985:nstate<=12'd986;
        12'd986:nstate<=12'd987;
        12'd987:nstate<=12'd988;
        12'd988:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd989;
                end
        12'd989:nstate<=12'd990;
        12'd990:nstate<=12'd991;
        12'd991:nstate<=12'd992;
        12'd992:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd993;
                end
        12'd993:nstate<=12'd994;
        12'd994:nstate<=12'd995;
        12'd995:nstate<=12'd996;
        12'd996:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd997;
                end
        12'd997:nstate<=12'd998;
        12'd998:nstate<=12'd999;
        12'd999:nstate<=12'd1000;
        12'd1000:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1001;
                end
        12'd1001:nstate<=12'd1002;
        12'd1002:nstate<=12'd1003;
        12'd1003:nstate<=12'd1004;
        12'd1004:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1005;
                end
        12'd1005:nstate<=12'd1006;
        12'd1006:nstate<=12'd1007;
        12'd1007:nstate<=12'd1008;
        12'd1008:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1009;
                end
        12'd1009:nstate<=12'd1010;
        12'd1010:nstate<=12'd1011;
        12'd1011:nstate<=12'd1012;
        12'd1012:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1013;
                end
        12'd1013:nstate<=12'd1014;
        12'd1014:nstate<=12'd1015;
        12'd1015:nstate<=12'd1016;
        12'd1016:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1017;
                end
        12'd1017:nstate<=12'd1018;
        12'd1018:nstate<=12'd1019;
        12'd1019:nstate<=12'd1020;
        12'd1020:
                        begin
                    if(indicator==1'd0)
                        nstate<=12'd1021;
                    else
                        nstate<=12'd1021;
                end
        default: nstate<=12'd1021;
        endcase
end


always@(*)
    begin
    case(pstate)
        12'd0:
            begin
                add_1<=8'd0;
                add_2<=8'd0;
                cin<=1'd0;
                en<=1'd0;
            end
        12'd1:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd0;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd2:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd3:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd4:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd5:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd1;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd6:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd7:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd8:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd9:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd2;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd10:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd11:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd12:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd13:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd3;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd14:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd15:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd16:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd17:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd4;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd18:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd19:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd20:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd21:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd5;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd22:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd23:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd24:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd25:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd6;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd26:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd27:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd28:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd29:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd7;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd30:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd31:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd32:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd33:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd8;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd34:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd35:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd36:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd37:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd9;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd38:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd39:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd40:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd41:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd10;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd42:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd43:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd44:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd45:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd11;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd46:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd47:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd48:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd49:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd12;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd50:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd51:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd52:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd53:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd13;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd54:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd55:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd56:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd57:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd14;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd58:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd59:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd60:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd61:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd15;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd62:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd63:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd64:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd65:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd16;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd66:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd67:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd68:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd69:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd17;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd70:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd71:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd72:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd73:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd18;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd74:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd75:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd76:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd77:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd19;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd78:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd79:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd80:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd81:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd20;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd82:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd83:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd84:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd85:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd21;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd86:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd87:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd88:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd89:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd22;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd90:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd91:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd92:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd93:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd23;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd94:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd95:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd96:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd97:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd24;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd98:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd99:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd100:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd101:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd25;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd102:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd103:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd104:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd105:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd26;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd106:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd107:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd108:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd109:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd27;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd110:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd111:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd112:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd113:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd28;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd114:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd115:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd116:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd117:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd29;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd118:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd119:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd120:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd121:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd30;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd122:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd123:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd124:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd125:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd31;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd126:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd127:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd128:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd129:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd32;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd130:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd131:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd132:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd133:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd33;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd134:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd135:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd136:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd137:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd34;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd138:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd139:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd140:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd141:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd35;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd142:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd143:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd144:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd145:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd36;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd146:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd147:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd148:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd149:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd37;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd150:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd151:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd152:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd153:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd38;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd154:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd155:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd156:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd157:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd39;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd158:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd159:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd160:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd161:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd40;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd162:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd163:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd164:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd165:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd41;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd166:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd167:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd168:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd169:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd42;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd170:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd171:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd172:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd173:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd43;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd174:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd175:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd176:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd177:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd44;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd178:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd179:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd180:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd181:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd45;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd182:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd183:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd184:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd185:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd46;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd186:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd187:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd188:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd189:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd47;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd190:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd191:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd192:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd193:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd48;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd194:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd195:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd196:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd197:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd49;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd198:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd199:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd200:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd201:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd50;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd202:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd203:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd204:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd205:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd51;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd206:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd207:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd208:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd209:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd52;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd210:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd211:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd212:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd213:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd53;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd214:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd215:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd216:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd217:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd54;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd218:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd219:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd220:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd221:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd55;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd222:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd223:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd224:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd225:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd56;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd226:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd227:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd228:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd229:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd57;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd230:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd231:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd232:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd233:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd58;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd234:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd235:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd236:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd237:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd59;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd238:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd239:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd240:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd241:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd60;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd242:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd243:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd244:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd245:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd61;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd246:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd247:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd248:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd249:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd62;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd250:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd251:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd252:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd253:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd63;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd254:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd255:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd256:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd257:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd64;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd258:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd259:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd260:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd261:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd65;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd262:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd263:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd264:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd265:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd66;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd266:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd267:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd268:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd269:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd67;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd270:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd271:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd272:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd273:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd68;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd274:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd275:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd276:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd277:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd69;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd278:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd279:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd280:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd281:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd70;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd282:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd283:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd284:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd285:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd71;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd286:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd287:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd288:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd289:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd72;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd290:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd291:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd292:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd293:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd73;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd294:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd295:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd296:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd297:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd74;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd298:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd299:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd300:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd301:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd75;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd302:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd303:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd304:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd305:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd76;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd306:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd307:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd308:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd309:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd77;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd310:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd311:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd312:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd313:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd78;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd314:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd315:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd316:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd317:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd79;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd318:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd319:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd320:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd321:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd80;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd322:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd323:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd324:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd325:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd81;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd326:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd327:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd328:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd329:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd82;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd330:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd331:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd332:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd333:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd83;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd334:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd335:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd336:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd337:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd84;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd338:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd339:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd340:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd341:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd85;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd342:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd343:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd344:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd345:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd86;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd346:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd347:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd348:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd349:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd87;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd350:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd351:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd352:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd353:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd88;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd354:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd355:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd356:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd357:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd89;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd358:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd359:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd360:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd361:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd90;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd362:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd363:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd364:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd365:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd91;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd366:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd367:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd368:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd369:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd92;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd370:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd371:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd372:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd373:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd93;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd374:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd375:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd376:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd377:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd94;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd378:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd379:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd380:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd381:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd95;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd382:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd383:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd384:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd385:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd96;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd386:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd387:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd388:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd389:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd97;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd390:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd391:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd392:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd393:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd98;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd394:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd395:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd396:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd397:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd99;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd398:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd399:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd400:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd401:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd100;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd402:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd403:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd404:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd405:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd101;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd406:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd407:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd408:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd409:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd102;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd410:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd411:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd412:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd413:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd103;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd414:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd415:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd416:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd417:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd104;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd418:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd419:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd420:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd421:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd105;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd422:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd423:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd424:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd425:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd106;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd426:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd427:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd428:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd429:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd107;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd430:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd431:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd432:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd433:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd108;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd434:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd435:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd436:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd437:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd109;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd438:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd439:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd440:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd441:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd110;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd442:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd443:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd444:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd445:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd111;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd446:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd447:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd448:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd449:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd112;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd450:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd451:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd452:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd453:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd113;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd454:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd455:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd456:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd457:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd114;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd458:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd459:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd460:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd461:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd115;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd462:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd463:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd464:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd465:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd116;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd466:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd467:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd468:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd469:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd117;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd470:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd471:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd472:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd473:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd118;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd474:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd475:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd476:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd477:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd119;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd478:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd479:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd480:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd481:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd120;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd482:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd483:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd484:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd485:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd121;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd486:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd487:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd488:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd489:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd122;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd490:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd491:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd492:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd493:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd123;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd494:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd495:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd496:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd497:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd124;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd498:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd499:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd500:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd501:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd125;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd502:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd503:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd504:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd505:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd126;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd506:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd507:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd508:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd509:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd127;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd510:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd511:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd512:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd513:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd128;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd514:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd515:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd516:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd517:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd129;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd518:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd519:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd520:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd521:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd130;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd522:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd523:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd524:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd525:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd131;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd526:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd527:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd528:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd529:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd132;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd530:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd531:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd532:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd533:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd133;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd534:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd535:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd536:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd537:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd134;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd538:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd539:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd540:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd541:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd135;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd542:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd543:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd544:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd545:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd136;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd546:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd547:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd548:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd549:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd137;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd550:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd551:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd552:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd553:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd138;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd554:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd555:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd556:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd557:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd139;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd558:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd559:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd560:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd561:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd140;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd562:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd563:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd564:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd565:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd141;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd566:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd567:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd568:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd569:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd142;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd570:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd571:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd572:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd573:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd143;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd574:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd575:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd576:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd577:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd144;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd578:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd579:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd580:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd581:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd145;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd582:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd583:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd584:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd585:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd146;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd586:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd587:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd588:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd589:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd147;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd590:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd591:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd592:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd593:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd148;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd594:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd595:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd596:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd597:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd149;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd598:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd599:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd600:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd601:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd150;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd602:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd603:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd604:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd605:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd151;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd606:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd607:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd608:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd609:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd152;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd610:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd611:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd612:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd613:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd153;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd614:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd615:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd616:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd617:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd154;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd618:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd619:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd620:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd621:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd155;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd622:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd623:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd624:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd625:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd156;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd626:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd627:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd628:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd629:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd157;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd630:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd631:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd632:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd633:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd158;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd634:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd635:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd636:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd637:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd159;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd638:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd639:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd640:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd641:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd160;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd642:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd643:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd644:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd645:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd161;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd646:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd647:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd648:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd649:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd162;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd650:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd651:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd652:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd653:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd163;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd654:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd655:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd656:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd657:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd164;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd658:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd659:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd660:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd661:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd165;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd662:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd663:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd664:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd665:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd166;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd666:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd667:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd668:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd669:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd167;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd670:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd671:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd672:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd673:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd168;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd674:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd675:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd676:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd677:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd169;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd678:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd679:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd680:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd681:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd170;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd682:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd683:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd684:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd685:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd171;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd686:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd687:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd688:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd689:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd172;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd690:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd691:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd692:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd693:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd173;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd694:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd695:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd696:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd697:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd174;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd698:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd699:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd700:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd701:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd175;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd702:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd703:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd704:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd705:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd176;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd706:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd707:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd708:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd709:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd177;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd710:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd711:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd712:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd713:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd178;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd714:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd715:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd716:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd717:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd179;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd718:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd719:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd720:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd721:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd180;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd722:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd723:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd724:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd725:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd181;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd726:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd727:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd728:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd729:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd182;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd730:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd731:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd732:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd733:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd183;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd734:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd735:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd736:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd737:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd184;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd738:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd739:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd740:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd741:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd185;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd742:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd743:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd744:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd745:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd186;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd746:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd747:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd748:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd749:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd187;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd750:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd751:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd752:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd753:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd188;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd754:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd755:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd756:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd757:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd189;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd758:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd759:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd760:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd761:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd190;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd762:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd763:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd764:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd765:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd191;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd766:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd767:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd768:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd769:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd192;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd770:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd771:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd772:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd773:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd193;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd774:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd775:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd776:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd777:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd194;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd778:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd779:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd780:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd781:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd195;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd782:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd783:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd784:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd785:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd196;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd786:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd787:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd788:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd789:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd197;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd790:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd791:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd792:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd793:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd198;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd794:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd795:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd796:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd797:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd199;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd798:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd799:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd800:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd801:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd200;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd802:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd803:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd804:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd805:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd201;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd806:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd807:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd808:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd809:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd202;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd810:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd811:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd812:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd813:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd203;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd814:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd815:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd816:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd817:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd204;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd818:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd819:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd820:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd821:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd205;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd822:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd823:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd824:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd825:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd206;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd826:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd827:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd828:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd829:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd207;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd830:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd831:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd832:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd833:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd208;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd834:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd835:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd836:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd837:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd209;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd838:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd839:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd840:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd841:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd210;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd842:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd843:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd844:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd845:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd211;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd846:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd847:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd848:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd849:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd212;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd850:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd851:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd852:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd853:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd213;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd854:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd855:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd856:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd857:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd214;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd858:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd859:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd860:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd861:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd215;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd862:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd863:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd864:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd865:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd216;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd866:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd867:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd868:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd869:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd217;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd870:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd871:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd872:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd873:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd218;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd874:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd875:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd876:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd877:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd219;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd878:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd879:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd880:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd881:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd220;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd882:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd883:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd884:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd885:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd221;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd886:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd887:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd888:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd889:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd222;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd890:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd891:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd892:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd893:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd223;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd894:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd895:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd896:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd897:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd224;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd898:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd899:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd900:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd901:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd225;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd902:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd903:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd904:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd905:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd226;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd906:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd907:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd908:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd909:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd227;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd910:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd911:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd912:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd913:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd228;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd914:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd915:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd916:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd917:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd229;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd918:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd919:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd920:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd921:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd230;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd922:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd923:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd924:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd925:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd231;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd926:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd927:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd928:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd929:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd232;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd930:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd931:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd932:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd933:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd233;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd934:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd935:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd936:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd937:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd234;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd938:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd939:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd940:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd941:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd235;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd942:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd943:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd944:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd945:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd236;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd946:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd947:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd948:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd949:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd237;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd950:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd951:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd952:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd953:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd238;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd954:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd955:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd956:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd957:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd239;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd958:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd959:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd960:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd961:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd240;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd962:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd963:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd964:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd965:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd241;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd966:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd967:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd968:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd969:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd242;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd970:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd971:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd972:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd973:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd243;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd974:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd975:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd976:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd977:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd244;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd978:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd979:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd980:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd981:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd245;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd982:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd983:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd984:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd985:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd246;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd986:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd987:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd988:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd989:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd247;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd990:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd991:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd992:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd993:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd248;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd994:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd995:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd996:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd997:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd249;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd998:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd999:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1000:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1001:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd250;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd1002:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1003:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1004:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1005:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd251;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd1006:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1007:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1008:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1009:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd252;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd1010:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1011:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1012:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1013:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd253;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd1014:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1015:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1016:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1017:
            begin
                add_1<=x_comp[7:0];
                add_2<=8'd254;
                cin<=1'd0;
                en<=1'd1;
            end
        12'd1018:
            begin
                add_1<=x_comp[15:8];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1019:
            begin
                add_1<=x_comp[23:16];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        12'd1020:
            begin
                add_1<=x_comp[31:24];
                add_2<=add_out;
                cin<=cout;
                en<=1'd1;
            end
        default:
            begin
                add_1<=add_1;
                add_2<=add_2;
                cin<=cin;
                en<=1'd0;
            end
        endcase
    end
 
endmodule
